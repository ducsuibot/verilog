module baitap_3_5_2(
	input wire [15:0] src1,
	input wire [15:0] src2,
	output [15:0] result
);
	assign result = src1 ^ src2; // Xor bit
endmodule