module baitap_3_5_1(
	input a, 
	input b,
	output out
);
	assign out = a&b;
endmodule