module baitap_3_5_7();
// mô phỏng các phép toán số học
  initial begin
    $display("5 + 10 = %d", 5 + 10);
    $display("5 - 10 = %d", 5 - 10);
    $display("10 - 5 = %d", 10 - 5);
    $display("10 * 5 = %d", 10 * 5);
    $display("10 / 5 = %d", 10 / 5);
    $display("10 / -5 = %d", 10 / -5);
    $display("10 %s 3 = %d", "%", 10 % 3);
    $display("+5 = %d", +5);
    $display("-5 = %d", -5);
    #10 $finish;
  end

endmodule